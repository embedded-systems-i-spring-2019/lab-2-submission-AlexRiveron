----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 03/07/2019 02:57:13 PM
-- Design Name: 
-- Module Name: my_alu - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use ieee.numeric_std.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity my_alu is
    Port ( A : in STD_LOGIC_VECTOR (3 downto 0);
           B : in STD_LOGIC_VECTOR (3 downto 0);
           opcode : in STD_LOGIC_VECTOR (3 downto 0);
           Y : out STD_LOGIC_VECTOR (3 downto 0));
end my_alu;

architecture Behavioral of my_alu is

begin
process (A,B,Opcode)
    begin
    
    case (opcode) is
    when "0000" => Y <= A+B;
    when "0001" => Y <= A-B;
    when "0010" => Y <= A+1;
    when "0011" => Y <= A-1;
    when "0100" => Y <= 0-A;
    when "0101" => if (A>B) then
                    Y <= "0001";
                 else
                    Y <= "0000";
                 end if;
    when "0110" => Y <= A(2 downto 0)&'0';
    when "0111" => Y <= '0' & A(3 downto 1);
    when "1000" => Y <= '1' & A(3 downto 1);
    when "1001" => Y <= not A;
    when "1010" => Y <= A and B;
    when "1011" => Y <= A or B;
    when "1100" => Y <= A xor B;
    when "1101" => Y <= A xnor B;
    when "1110" => Y <= A nand B;
    when "1111" => Y <= A nor B;
    end case;
end process;

end Behavioral;
